*bp_4stage.cir -- 4-stage bandpass filter
* 13 ideal opamps

R1 1 2 1
R2 13 3 1
R3 2 0 1
R4 3 4 1
E1 4 0 2 3 10G

R5 4 5 1
R6 5 6 1
C6 5 6 100u
E2 6 0 0 5 10G

R7 6 7 1
C8 7 8 100u
E3 8 0 0 7 10G

R9 8 3 1

R10 6 9 1
R11 20 10 1
R12 9 0 1
R13 10 11 1
E4 11 0 9 10 10G

R14 11 12 1
R15 12 13 1
C15 12 13 100u
E5 13 0 0 12 10G

R16 13 14 1
C17 14 15 100u
E6 15 0 0 14 10G

R18 15 10 1

R19 13 16 1
R20 17 27 1
R21 16 0 1
R22 17 18 1
E7 18 0 16 17 10G

R23 18 19 1
R24 19 20 1
C24 19 20 100u
E8 20 0 0 19 10G

R25 20 21 1
C26 21 22 100u
E9 22 0 0 21 10G

R27 22 17 1

R28 20 23 1
R29 32 24 1
R30 23 0  1
R31 24 25 1
E10 25 0 23 24 10G

R32 25 26 1
R33 26 27 1
C33 26 27 100u
E11 27 0 0 26 10G

R34 27 28 1
C35 28 29 100u
E12 29 0 0 28 10G

R36 29 24 1

R37 27 30 1
R38 0 31 1 
R39 0 30 1
R40 31 32 1
E13 32 0 30 31 10G

Vin 1 0 1
.ac 32 0 dec 2 1 10meg
.end

